000000000192   ���� �������� ������ ����� ����                                                                                                                                                                                                                                19                                                                                                                                                                                                                                                             
Fault5.wav                                                                                                                                                                                                                                                     000000000208   $�������� ���������� ����� ����� ����                                                                                                                                                                                                                           20                                                                                                                                                                                                                                                             Fault122.wav                                                                                                                                                                                                                                                   000000000215   ���� ���������� ����������                                                                                                                                                                                                                                     21                                                                                                                                                                                                                                                             Fault11.wav                                                                                                                                                                                                                                                    000000000222   ������� � ���� � �������                                                                                                                                                                                                                                       22                                                                                                                                                                                                                                                             Fault123.wav                                                                                                                                                                                                                                                   000000000185   $������������� ��� �������� ���������                                                                                                                                                                                                                           18                                                                                                                                                                                                                                                             Fault18.wav                                                                                                                                                                                                                                                    000000000239   ���� �� ��� ���� ����������                                                                                                                                                                                                                                    23                                                                                                                                                                                                                                                             
Fault6.wav                                                                                                                                                                                                                                                     000000000253   
���� �����                                                                                                                                                                                                                                                     25                                                                                                                                                                                                                                                             Fault125.wav                                                                                                                                                                                                                                                   000000000260   ���� ����������� ������ �����                                                                                                                                                                                                                                  26                                                                                                                                                                                                                                                             Fault126.wav                                                                                                                                                                                                                                                   000000000277   ������������� � ���� �����                                                                                                                                                                                                                                     27                                                                                                                                                                                                                                                             Fault127.wav                                                                                                                                                                                                                                                   000000000062   �� �������� � ����� ������                                                                                                                                                                                                                                     6                                                                                                                                                                                                                                                              Fault17.wav                                                                                                                                                                                                                                                    000000000130   �������� ����� ����������                                                                                                                                                                                                                                      13                                                                                                                                                                                                                                                             Fault118.wav                                                                                                                                                                                                                                                   000000000031   $������ �������� ����, ���� ��� �����                                                                                                                                                                                                                           3                                                                                                                                                                                                                                                              Fault112.wav                                                                                                                                                                                                                                                   000000000048   %������ �������� ����, ���� ��� ������                                                                                                                                                                                                                          4                                                                                                                                                                                                                                                              Fault113.wav                                                                                                                                                                                                                                                   000000000017   ������������� ��� ������                                                                                                                                                                                                                                       1                                                                                                                                                                                                                                                              Fault111.wav                                                                                                                                                                                                                                                   000000000055   �������������� ������                                                                                                                                                                                                                                          5                                                                                                                                                                                                                                                              Fault114.wav                                                                                                                                                                                                                                                   000000000178   ,��������� ����������� ����������� ����������                                                                                                                                                                                                                   17                                                                                                                                                                                                                                                             Fault14.wav                                                                                                                                                                                                                                                    000000000024   ����������� ���� ��� ������                                                                                                                                                                                                                                    2                                                                                                                                                                                                                                                              Fault10.wav                                                                                                                                                                                                                                                    000000000116   �������� ��������� ����������                                                                                                                                                                                                                                  11                                                                                                                                                                                                                                                             Fault116.wav                                                                                                                                                                                                                                                   000000000093   �� �������� �����                                                                                                                                                                                                                                              9                                                                                                                                                                                                                                                              Fault16.wav                                                                                                                                                                                                                                                    000000000123   ��� ���������� ���������� �����                                                                                                                                                                                                                                12                                                                                                                                                                                                                                                             Fault117.wav                                                                                                                                                                                                                                                   000000000086   �� �������� � ������ ������                                                                                                                                                                                                                                    8                                                                                                                                                                                                                                                              Fault13.wav                                                                                                                                                                                                                                                    000000000109   $�������� � ������ ������� ����������                                                                                                                                                                                                                           10                                                                                                                                                                                                                                                             Fault115.wav                                                                                                                                                                                                                                                   000000000161   �� ���������� ����������� �����                                                                                                                                                                                                                                16                                                                                                                                                                                                                                                             Fault121.wav                                                                                                                                                                                                                                                   000000000147   ����� ���������� ��� ����������                                                                                                                                                                                                                                14                                                                                                                                                                                                                                                             Fault119.wav                                                                                                                                                                                                                                                   000000000079   �� �������� � ������ ������                                                                                                                                                                                                                                    7                                                                                                                                                                                                                                                              
Fault7.wav                                                                                                                                                                                                                                                     000000000246   ������ ��� ��� ����������                                                                                                                                                                                                                                      24                                                                                                                                                                                                                                                             Fault124.wav                                                                                                                                                                                                                                                   000000000154   "��������� ��������� � ���� �������                                                                                                                                                                                                                             15                                                                                                                                                                                                                                                             Fault120.wav                                                                                                                                                                                                                                                   